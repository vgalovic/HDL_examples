library IEEE;
  use IEEE.STD_LOGIC_1164.ALL;
  use IEEE.NUMERIC_STD.ALL;
  use IEEE.MATH_REAL.ALL;

entity mod_100_counter_down is
    Generic (
        M : integer := 100;
        WIDTH : integer := integer(ceil(log2(real(100))))
    );
    Port (
        clk : in STD_LOGIC;
        ce, en : in STD_LOGIC;
        load : in STD_LOGIC;
        counter_value: in  STD_LOGIC_VECTOR(WIDTH -1 downto 0);
        q : out STD_LOGIC_VECTOR (WIDTH - 1 downto 0)
    );
end mod_100_counter_down;

architecture Behavioral of mod_100_counter_down is
    subtype cnt_range_t is integer range 0 to M - 1;
    signal count_s : cnt_range_t := M - 1;

begin
    cnt: process(clk, ce, en, load, count_s, counter_value)
    begin
        if rising_edge(clk) then
            if ce = '1' then
                if load = '1' then
                    if counter_value <  std_logic_vector(to_unsigned(M, WIDTH)) then
                        count_s <= to_integer(unsigned(counter_value(WIDTH - 1 downto 0)));
                    end if;
                elsif en = '1' then
                    if count_s = 0 then
                        count_s <= M - 1;
                    else
                        count_s <= count_s - 1;
                    end if;
                end if;
            end if;
        end if;
    end process cnt;

    q <= std_logic_vector(to_unsigned(count_s, WIDTH));

end Behavioral;
